`timescale 1ns/1ns

module fft_256_tb (
    output logic clk
);

localparam WIDTH = 12;  // time-domain sample width
localparam N = 256;     // FFT points

logic rst, start, done;

logic [WIDTH-1:0] time_samples [0:N-1] = '{
-32, -185, -128, -178, 99, -125, 160, 63, -38, -105, -125, 13, -153, 119, 87, 18, -76, -84, 93, -33, -5, -98, 60, 163, -149, 159, -162, -167, -142, 180, 55, 123, 125, -112, -4, 102, 151, 11, -79, -169, -120, -148, 38, -150, -68, 18, 119, 7, -151, 95, -64, 71, 33, 192, 47, 48, 173, -127, -15, 161, 166, 52, -117, -104, -157, 88, -174, 192, -124, 54, -62, 96, -166, 116, -63, 46, 126, -114, -181, -144, 185, 124, -32, -119, -139, -75, -103, 143, 99, 108, 29, 18, 24, -184, 111, -77, -51, -157, 8, 126, 2, -141, 73, -57, -42, -174, 95, 119, 39, -52, -13, -23, 156, 50, 55, -173, -200, -138, 45, -108, 92, -137, -125, -90, -150, 1, -65, 49, 138, 185, 7, 19, 38, 24, -151, 96, 164, -154, 129, -122, -90, -105, 88, 175, 72, -142, -179, 34, -9, 11, 148, -149, -103, -192, -93, -114, -112, 167, -61, 57, -3, 115, -137, -65, 136, 161, 148, 7, -78, -55, 113, 90, 98, -152, -164, -178, -181, -105, -155, 128, 93, -191, -51, 42, 139, 146, -164, 96, 158, -181, -16, 192, 180, 6, 173, -151, -149, -85, -5, -121, 186, 78, 61, -67, 10, 157, 149, -60, 20, 190, -87, -156, -195, -3, 108, 176, 118, 139, 159, -99, -47, -75, -164, -57, 13, 74, 78, -107, 70, -136, -113, 89, 158, -129, -104, -118, -121, 146, 8, 62, 53, 190, -15, 41, 141, -95, -36, 33, -137, -96, 11, -196, 110, 52, -78, 55
};

logic [WIDTH:0] freq_real [0:N-1];
logic [WIDTH:0] freq_imag [0:N-1];
logic [WIDTH+1:0] freq_mag [0:N-1];

fft_256 #(.WIDTH(WIDTH)) DUT (
    .clk(clk),
    .rst(rst),
    .start(start),
    .done(done),
    .time_samples(time_samples),
    .freq_real(freq_real),
    .freq_imag(freq_imag)
);

mag_est #(.WIDTH(WIDTH)) EST (
    .real_in(freq_real),
    .imag_in(freq_imag),
    .magnitude(freq_mag)
);

initial begin
    clk <= 0;
    rst <= 1;
    start <= 0;

    #10 rst <= 0;
    start <= 1;
	 #10 start <= 0;

    #70 rst <= 1;
	 #10 rst <= 0;
	 #10 start <= 1;
	 #10 start <= 0;
	 
	 #80 $stop;
end

always begin
    #5 clk = ~clk;
end

endmodule