`timescale 1ns/1ns

module fft_256_tb (
    output logic clk
);

localparam WIDTH = 20;  // computation bit width
localparam N = 256;     // FFT points

logic [WIDTH-1:0] time_samples [0:N-1] = '{
    1061, 235, 3980, 1096, 3839, 905, 2763, 3717, 2895, 960, 144, 129, 4044, 3655, 2797, 2556, 3462, 3353, 1202, 1300, 1278, 357, 2962, 2516, 2955, 252, 3562, 668, 3997, 2446, 562, 2628, 3287, 4055, 3049, 753, 1527, 3550, 1888, 1110, 2189, 2025, 3465, 1031, 319, 2877, 3606, 1337, 2561, 1920, 316, 2257, 1288, 728, 3725, 2675, 431, 4074, 633, 2504, 542, 1095, 1411, 1478, 3989, 3633, 1337, 515, 3012, 2840, 497, 3115, 1612, 3098, 1844, 1360, 2669, 883, 1321, 3538, 15, 3136, 2244, 25, 3439, 3810, 1495, 1927, 1306, 3737, 1640, 1046, 1801, 3779, 3047, 1150, 1303, 3453, 3428, 155, 2981, 313, 2643, 3238, 648, 1312, 3490, 3850, 3351, 1679, 2799, 3159, 3865, 4039, 243, 1372, 2634, 1214, 3374, 928, 1752, 1175, 695, 1345, 1393, 1869, 1795, 2944, 4088, 1277, 461, 1798, 564, 469, 1478, 1538, 1612, 4059, 2197, 715, 2311, 2125, 2760, 1099, 3404, 1067, 532, 3614, 1572, 871, 1799, 3885, 964, 2617, 3824, 3580, 2258, 96, 269, 3082, 2327, 3964, 2897, 1927, 889, 152, 1738, 3548, 3732, 2464, 3212, 3265, 606, 3644, 489, 152, 3410, 883, 865, 2178, 3564, 1756, 2663, 1890, 266, 3766, 1888, 2537, 1874, 2518, 3270, 2754, 327, 4071, 2224, 1590, 3087, 2949, 1425, 2218, 20, 2678, 1968, 2326, 2533, 3981, 2033, 2674, 609, 1717, 1876, 3082, 3168, 183, 2365, 3640, 3801, 405, 3303, 3168, 505, 4051, 1049, 1521, 910, 2189, 3284, 3700, 811, 3718, 1741, 696, 1979, 2959, 1560, 1019, 3209, 450, 2247, 3893, 3397, 2468, 869, 2808, 2069, 3368, 77, 2267, 2737, 2417, 1327, 1485, 3496, 1486, 1581, 1879
};

logic rst, start;
logic done, done_old;

logic [WIDTH:0] freq_mag [0:N-1];
logic [WIDTH:0] freq_mag_old [0:N-1];

fft_256 #(.WIDTH(WIDTH)) DUT (
    .clk(clk),
    .rst(rst),
    .start(start),
    .done(done),
    .time_samples(time_samples),
    .freq_mag(freq_mag)
);

// fft_256_old #(.WIDTH(WIDTH)) OLD (
//     .clk(clk),
//     .rst(rst),
//     .start(start),
//     .done(done_old),
//     .time_samples(time_samples),
//     .freq_mag(freq_mag_old)
// );

// mag_est #(.WIDTH(WIDTH)) EST_OLD (
//     .real_in(freq_real_old),
//     .imag_in(freq_imag_old),
//     .magnitude(freq_mag_old)
// );

initial begin
    clk <= 0;
    rst <= 1;
    start <= 0;

    #10 rst <= 0;
    start <= 1;
	#10 start <= 0;

    #1000 rst <= 1;
	#10 rst <= 0;
	#10 start <= 1;
	#10 start <= 0;
	
	#80 $stop;
end

always begin
    #5 clk = ~clk;
end

endmodule