module fft_256 #(
    parameter WIDTH = 18,
    parameter USED_SAMPLES = 256, // number of frequency bins to output
    parameter N = 256  // must be power of 4
) (
    input clk,
    input rst,
    input start,
    output done,

    input [WIDTH-1:0] time_samples [0:N-1],
    output logic [WIDTH:0] freq_mag [0:USED_SAMPLES-1]
);

/*
    256-point decimation-in-time FFT using radix-4 butterfly units. 
    64 butterfly units are needed, but due to device (Intel MAX10 10M50DAF484C7G) limitations, we can only instantiate 16 at a time. 
    each stage is split into four sub-stages to perform computations in parallel. 
    12b twiddle factor (plus sign bit) is necessary to retain uniqueness of finest granularity twiddle factors.
    increased width yields higher accuracy at the cost of more resources.
    this module assumes a 12b input bus of time-domain data, and outputs a 18b bus of approximated complex frequency magnitudes. 

    TODO: look into loading ROM for twiddle factors? not sure if read latency will be an issue, currently stored in logic array

    handy resources for 4-radix FFT implementations: 
        https://www.ti.com/lit/an/spra152/spra152.pdf 
        https://www.cmlab.csie.ntu.edu.tw/cml/dsp/training/coding/transform/fft.html
        https://thescipub.com/abstract/ajassp.2007.570.575 
        https://www.worldscientific.com/doi/abs/10.1142/S021812661240018X
*/

localparam N_BFLY = (N+3)/4;
localparam N_INST = 4;
localparam N_LOG2 = $clog2(N);
localparam N_STAGES = N_LOG2/2;
localparam FULL_WIDTH = WIDTH*2;

// inputs to instantiated butterfly units
logic [0:N_INST-1] [FULL_WIDTH-1:0] a;
logic [0:N_INST-1] [FULL_WIDTH-1:0] b;
logic [0:N_INST-1] [FULL_WIDTH-1:0] c;
logic [0:N_INST-1] [FULL_WIDTH-1:0] d;
logic [0:N_INST-1] [FULL_WIDTH-1:0] w0;
logic [0:N_INST-1] [FULL_WIDTH-1:0] w1;
logic [0:N_INST-1] [FULL_WIDTH-1:0] w2;
logic [0:N_INST-1] [FULL_WIDTH-1:0] w3;

// outputs of instantiated butterfly units
logic [0:N_INST-1] [FULL_WIDTH-1:0] out_d [0:3];

// outputs of butterfly units 0:N_BFLY-1 from previous stage
logic [0:N_BFLY-1] [FULL_WIDTH-1:0] out_temp [0:3]; 
logic [0:N_BFLY-1] [FULL_WIDTH-1:0] out [0:3];

// twiddle factors for 256-point FFT, generated by gen_twiddle.py
logic [0:189] [FULL_WIDTH-1:0] w_256 = '{
        { 18'd131071,    18'd0},        // W0
        { 18'd131032,   -18'd3216},     // W1
        { 18'd130914,   -18'd6431},     // W2
        { 18'd130716,   -18'd9642},     // W3
        { 18'd130440,   -18'd12847},    // W4
        { 18'd130086,   -18'd16044},    // W5
        { 18'd129653,   -18'd19232},    // W6
        { 18'd129142,   -18'd22408},    // W7
        { 18'd128553,   -18'd25570},    // W8
        { 18'd127887,   -18'd28718},    // W9
        { 18'd127143,   -18'd31847},    // W10
        { 18'd126324,   -18'd34958},    // W11
        { 18'd125428,   -18'd38048},    // W12
        { 18'd124456,   -18'd41114},    // W13
        { 18'd123410,   -18'd44156},    // W14
        { 18'd122289,   -18'd47172},    // W15
        { 18'd121094,   -18'd50159},    // W16
        { 18'd119827,   -18'd53115},    // W17
        { 18'd118487,   -18'd56040},    // W18
        { 18'd117076,   -18'd58931},    // W19
        { 18'd115595,   -18'd61786},    // W20
        { 18'd114044,   -18'd64605},    // W21
        { 18'd112424,   -18'd67384},    // W22
        { 18'd110736,   -18'd70123},    // W23
        { 18'd108982,   -18'd72819},    // W24
        { 18'd107162,   -18'd75472},    // W25
        { 18'd105278,   -18'd78079},    // W26
        { 18'd103330,   -18'd80639},    // W27
        { 18'd101320,   -18'd83151},    // W28
        { 18'd99248,    -18'd85612},    // W29
        { 18'd97117,    -18'd88022},    // W30
        { 18'd94928,    -18'd90379},    // W31
        { 18'd92681,    -18'd92681},    // W32
        { 18'd90379,    -18'd94928},    // W33
        { 18'd88022,    -18'd97117},    // W34
        { 18'd85612,    -18'd99248},    // W35
        { 18'd83151,    -18'd101320},   // W36
        { 18'd80639,    -18'd103330},   // W37
        { 18'd78079,    -18'd105278},   // W38
        { 18'd75472,    -18'd107162},   // W39
        { 18'd72819,    -18'd108982},   // W40
        { 18'd70123,    -18'd110736},   // W41
        { 18'd67384,    -18'd112424},   // W42
        { 18'd64605,    -18'd114044},   // W43
        { 18'd61786,    -18'd115595},   // W44
        { 18'd58931,    -18'd117076},   // W45
        { 18'd56040,    -18'd118487},   // W46
        { 18'd53115,    -18'd119827},   // W47
        { 18'd50159,    -18'd121094},   // W48
        { 18'd47172,    -18'd122289},   // W49
        { 18'd44156,    -18'd123410},   // W50
        { 18'd41114,    -18'd124456},   // W51
        { 18'd38048,    -18'd125428},   // W52
        { 18'd34958,    -18'd126324},   // W53
        { 18'd31847,    -18'd127143},   // W54
        { 18'd28718,    -18'd127887},   // W55
        { 18'd25570,    -18'd128553},   // W56
        { 18'd22408,    -18'd129142},   // W57
        { 18'd19232,    -18'd129653},   // W58
        { 18'd16044,    -18'd130086},   // W59
        { 18'd12847,    -18'd130440},   // W60
        { 18'd9642,     -18'd130716},   // W61
        { 18'd6431,     -18'd130914},   // W62
        { 18'd3216,     -18'd131032},   // W63
        { 18'd0,        -18'd131072},   // W64
        {-18'd3216,     -18'd131032},   // W65
        {-18'd6431,     -18'd130914},   // W66
        {-18'd9642,     -18'd130716},   // W67
        {-18'd12847,    -18'd130440},   // W68
        {-18'd16044,    -18'd130086},   // W69
        {-18'd19232,    -18'd129653},   // W70
        {-18'd22408,    -18'd129142},   // W71
        {-18'd25570,    -18'd128553},   // W72
        {-18'd28718,    -18'd127887},   // W73
        {-18'd31847,    -18'd127143},   // W74
        {-18'd34958,    -18'd126324},   // W75
        {-18'd38048,    -18'd125428},   // W76
        {-18'd41114,    -18'd124456},   // W77
        {-18'd44156,    -18'd123410},   // W78
        {-18'd47172,    -18'd122289},   // W79
        {-18'd50159,    -18'd121094},   // W80
        {-18'd53115,    -18'd119827},   // W81
        {-18'd56040,    -18'd118487},   // W82
        {-18'd58931,    -18'd117076},   // W83
        {-18'd61786,    -18'd115595},   // W84
        {-18'd64605,    -18'd114044},   // W85
        {-18'd67384,    -18'd112424},   // W86
        {-18'd70123,    -18'd110736},   // W87
        {-18'd72819,    -18'd108982},   // W88
        {-18'd75472,    -18'd107162},   // W89
        {-18'd78079,    -18'd105278},   // W90
        {-18'd80639,    -18'd103330},   // W91
        {-18'd83151,    -18'd101320},   // W92
        {-18'd85612,    -18'd99248},    // W93
        {-18'd88022,    -18'd97117},    // W94
        {-18'd90379,    -18'd94928},    // W95
        {-18'd92681,    -18'd92681},    // W96
        {-18'd94928,    -18'd90379},    // W97
        {-18'd97117,    -18'd88022},    // W98
        {-18'd99248,    -18'd85612},    // W99
        {-18'd101320,   -18'd83151},    // W100
        {-18'd103330,   -18'd80639},    // W101
        {-18'd105278,   -18'd78079},    // W102
        {-18'd107162,   -18'd75472},    // W103
        {-18'd108982,   -18'd72819},    // W104
        {-18'd110736,   -18'd70123},    // W105
        {-18'd112424,   -18'd67384},    // W106
        {-18'd114044,   -18'd64605},    // W107
        {-18'd115595,   -18'd61786},    // W108
        {-18'd117076,   -18'd58931},    // W109
        {-18'd118487,   -18'd56040},    // W110
        {-18'd119827,   -18'd53115},    // W111
        {-18'd121094,   -18'd50159},    // W112
        {-18'd122289,   -18'd47172},    // W113
        {-18'd123410,   -18'd44156},    // W114
        {-18'd124456,   -18'd41114},    // W115
        {-18'd125428,   -18'd38048},    // W116
        {-18'd126324,   -18'd34958},    // W117
        {-18'd127143,   -18'd31847},    // W118
        {-18'd127887,   -18'd28718},    // W119
        {-18'd128553,   -18'd25570},    // W120
        {-18'd129142,   -18'd22408},    // W121
        {-18'd129653,   -18'd19232},    // W122
        {-18'd130086,   -18'd16044},    // W123
        {-18'd130440,   -18'd12847},    // W124
        {-18'd130716,   -18'd9642},     // W125
        {-18'd130914,   -18'd6431},     // W126
        {-18'd131032,   -18'd3216},     // W127
        {-18'd131072,    18'd0},        // W128
        {-18'd131032,    18'd3216},     // W129
        {-18'd130914,    18'd6431},     // W130
        {-18'd130716,    18'd9642},     // W131
        {-18'd130440,    18'd12847},    // W132
        {-18'd130086,    18'd16044},    // W133
        {-18'd129653,    18'd19232},    // W134
        {-18'd129142,    18'd22408},    // W135
        {-18'd128553,    18'd25570},    // W136
        {-18'd127887,    18'd28718},    // W137
        {-18'd127143,    18'd31847},    // W138
        {-18'd126324,    18'd34958},    // W139
        {-18'd125428,    18'd38048},    // W140
        {-18'd124456,    18'd41114},    // W141
        {-18'd123410,    18'd44156},    // W142
        {-18'd122289,    18'd47172},    // W143
        {-18'd121094,    18'd50159},    // W144
        {-18'd119827,    18'd53115},    // W145
        {-18'd118487,    18'd56040},    // W146
        {-18'd117076,    18'd58931},    // W147
        {-18'd115595,    18'd61786},    // W148
        {-18'd114044,    18'd64605},    // W149
        {-18'd112424,    18'd67384},    // W150
        {-18'd110736,    18'd70123},    // W151
        {-18'd108982,    18'd72819},    // W152
        {-18'd107162,    18'd75472},    // W153
        {-18'd105278,    18'd78079},    // W154
        {-18'd103330,    18'd80639},    // W155
        {-18'd101320,    18'd83151},    // W156
        {-18'd99248,     18'd85612},    // W157
        {-18'd97117,     18'd88022},    // W158
        {-18'd94928,     18'd90379},    // W159
        {-18'd92681,     18'd92681},    // W160
        {-18'd90379,     18'd94928},    // W161
        {-18'd88022,     18'd97117},    // W162
        {-18'd85612,     18'd99248},    // W163
        {-18'd83151,     18'd101320},   // W164
        {-18'd80639,     18'd103330},   // W165
        {-18'd78079,     18'd105278},   // W166
        {-18'd75472,     18'd107162},   // W167
        {-18'd72819,     18'd108982},   // W168
        {-18'd70123,     18'd110736},   // W169
        {-18'd67384,     18'd112424},   // W170
        {-18'd64605,     18'd114044},   // W171
        {-18'd61786,     18'd115595},   // W172
        {-18'd58931,     18'd117076},   // W173
        {-18'd56040,     18'd118487},   // W174
        {-18'd53115,     18'd119827},   // W175
        {-18'd50159,     18'd121094},   // W176
        {-18'd47172,     18'd122289},   // W177
        {-18'd44156,     18'd123410},   // W178
        {-18'd41114,     18'd124456},   // W179
        {-18'd38048,     18'd125428},   // W180
        {-18'd34958,     18'd126324},   // W181
        {-18'd31847,     18'd127143},   // W182
        {-18'd28718,     18'd127887},   // W183
        {-18'd25570,     18'd128553},   // W184
        {-18'd22408,     18'd129142},   // W185
        {-18'd19232,     18'd129653},   // W186
        {-18'd16044,     18'd130086},   // W187
        {-18'd12847,     18'd130440},   // W188
        {-18'd9642,      18'd130716}    // W189
};

// frequency output magnitude estimation
logic [WIDTH-1:0] freq_real [0:N-1];
logic [WIDTH-1:0] freq_imag [0:N-1];
mag_est #(.WIDTH(WIDTH), .N(USED_SAMPLES)) MAG ( 
	.real_in(freq_real[0:USED_SAMPLES-1]), 
	.imag_in(freq_imag[0:USED_SAMPLES-1]), 
	.magnitude(freq_mag[0:USED_SAMPLES-1])
);

typedef enum logic [2:0] {SET, STAGE1, STAGE2, STAGE3, STAGE4, DONE} state_t;
state_t state, state_d;
logic [3:0] counter;
logic [1:0] substage;
logic [1:0] subsubstage;
assign substage = counter[3:2];
assign subsubstage = counter[1:0];

logic [1:0] done_sr;
assign done = (state == DONE);

// INSTANTIATE RADIX4 BFLY UNITS
genvar i;
generate 
    for (i = 0; i < N_INST; i++) begin : gen_BFLY
        butterfly_4 #(.FULL_WIDTH(FULL_WIDTH)) butterfly (
            .a(a[i]),
            .b(b[i]),
            .c(c[i]),
            .d(d[i]),
            .w0(w0[i]),
            .w1(w1[i]),
            .w2(w2[i]),
            .w3(w3[i]),
            .out0(out_d[0][i]),
            .out1(out_d[1][i]),
            .out2(out_d[2][i]),
            .out3(out_d[3][i])
        );
    end
endgenerate

always_ff @(posedge clk) begin
    if (rst) begin
        done_sr <= 2'b0;
        state <= SET;
        counter <= 2'b00;
    end else begin
        done_sr <= {(state_d == DONE), done_sr[1]};
        state <= state_d;
        counter <= counter + ((state == SET) ? 1'b0 : 1'b1);
    end

    // update out using temp array
    if (state != state_d) begin
        out <= out_temp;
    end
end

// update temp array of stage outputs with substaged butterfly outputs
always_ff @(negedge clk) begin

    case (counter)
    4'h0: begin
        out_temp[0][0:3] <= out_d[0];
        out_temp[1][0:3] <= out_d[1];
        out_temp[2][0:3] <= out_d[2];
        out_temp[3][0:3] <= out_d[3];
    end
    4'h1: begin
        out_temp[0][4:7] <= out_d[0];
        out_temp[1][4:7] <= out_d[1];
        out_temp[2][4:7] <= out_d[2];
        out_temp[3][4:7] <= out_d[3];
    end
    4'h2: begin
        out_temp[0][8:11] <= out_d[0];
        out_temp[1][8:11] <= out_d[1];
        out_temp[2][8:11] <= out_d[2];
        out_temp[3][8:11] <= out_d[3];
    end
    4'h3: begin
        out_temp[0][12:15] <= out_d[0];
        out_temp[1][12:15] <= out_d[1];
        out_temp[2][12:15] <= out_d[2];
        out_temp[3][12:15] <= out_d[3];
    end
    4'h4: begin
        out_temp[0][16:19] <= out_d[0];
        out_temp[1][16:19] <= out_d[1];
        out_temp[2][16:19] <= out_d[2];
        out_temp[3][16:19] <= out_d[3];
    end
    4'h5: begin
        out_temp[0][20:23] <= out_d[0];
        out_temp[1][20:23] <= out_d[1];
        out_temp[2][20:23] <= out_d[2];
        out_temp[3][20:23] <= out_d[3];
    end
    4'h6: begin
        out_temp[0][24:27] <= out_d[0];
        out_temp[1][24:27] <= out_d[1];
        out_temp[2][24:27] <= out_d[2];
        out_temp[3][24:27] <= out_d[3];
    end
    4'h7: begin
        out_temp[0][28:31] <= out_d[0];
        out_temp[1][28:31] <= out_d[1];
        out_temp[2][28:31] <= out_d[2];
        out_temp[3][28:31] <= out_d[3];
    end
    4'h8: begin
        out_temp[0][32:35] <= out_d[0];
        out_temp[1][32:35] <= out_d[1];
        out_temp[2][32:35] <= out_d[2];
        out_temp[3][32:35] <= out_d[3];
    end
    4'h9: begin
        out_temp[0][36:39] <= out_d[0];
        out_temp[1][36:39] <= out_d[1];
        out_temp[2][36:39] <= out_d[2];
        out_temp[3][36:39] <= out_d[3];
    end
    4'ha: begin
        out_temp[0][40:43] <= out_d[0];
        out_temp[1][40:43] <= out_d[1];
        out_temp[2][40:43] <= out_d[2];
        out_temp[3][40:43] <= out_d[3];
    end
    4'hb: begin
        out_temp[0][44:47] <= out_d[0];
        out_temp[1][44:47] <= out_d[1];
        out_temp[2][44:47] <= out_d[2];
        out_temp[3][44:47] <= out_d[3];
    end
    4'hc: begin
        out_temp[0][48:51] <= out_d[0];
        out_temp[1][48:51] <= out_d[1];
        out_temp[2][48:51] <= out_d[2];
        out_temp[3][48:51] <= out_d[3];
    end
    4'hd: begin
        out_temp[0][52:55] <= out_d[0];
        out_temp[1][52:55] <= out_d[1];
        out_temp[2][52:55] <= out_d[2];
        out_temp[3][52:55] <= out_d[3];
    end
    4'he: begin
        out_temp[0][56:59] <= out_d[0];
        out_temp[1][56:59] <= out_d[1];
        out_temp[2][56:59] <= out_d[2];
        out_temp[3][56:59] <= out_d[3];
    end
    4'hf: begin
        out_temp[0][60:63] <= out_d[0];
        out_temp[1][60:63] <= out_d[1];
        out_temp[2][60:63] <= out_d[2];
        out_temp[3][60:63] <= out_d[3];
    end
    default: begin
        out_temp[0] <= 1'b0;
        out_temp[1] <= 1'b0;
        out_temp[2] <= 1'b0;
        out_temp[3] <= 1'b0;
    end
    endcase
end

// state machine for butterfly unit inputs
always_comb begin
    case (state) 
    SET: begin
        for (int i = 0; i < N_INST; i++) begin
            a[i] = 1'b0;
            b[i] = 1'b0;
            c[i] = 1'b0;
            d[i] = 1'b0;
            w0[i]= 1'b0;
            w1[i]= 1'b0;
            w2[i]= 1'b0;
            w3[i]= 1'b0;
        end
    end

    STAGE1: begin   
        for (int i = 0; i < N_INST; i++) begin
            a[i][FULL_WIDTH-1:WIDTH] = 1'd0 + time_samples[i+N_BFLY*0+substage*16+subsubstage*4];
            b[i][FULL_WIDTH-1:WIDTH] = 1'd0 + time_samples[i+N_BFLY*1+substage*16+subsubstage*4];
            c[i][FULL_WIDTH-1:WIDTH] = 1'd0 + time_samples[i+N_BFLY*2+substage*16+subsubstage*4];
            d[i][FULL_WIDTH-1:WIDTH] = 1'd0 + time_samples[i+N_BFLY*3+substage*16+subsubstage*4];
            a[i][WIDTH-1:0] = 1'b0;
            b[i][WIDTH-1:0] = 1'b0;
            c[i][WIDTH-1:0] = 1'b0;
            d[i][WIDTH-1:0] = 1'b0;
            w0[i] = w_256[0];
            w1[i] = w_256[0];
            w2[i] = w_256[0];
            w3[i] = w_256[0];
        end
    end

    STAGE2: begin
        // for (int i = 0; i < 4; i++) begin
        //     for (int j = 0; j < 16; j++) begin
        //         a[i*16+j] = out[i][j+0*16];
        //         b[i*16+j] = out[i][j+1*16];
        //         c[i*16+j] = out[i][j+2*16];
        //         d[i*16+j] = out[i][j+3*16];
        //         w0[i*16+j]= w_256[i*(j+0*16)];
        //         w1[i*16+j]= w_256[i*(j+1*16)];
        //         w2[i*16+j]= w_256[i*(j+2*16)];
        //         w3[i*16+j]= w_256[i*(j+3*16)];
        //     end
        // end
        for (int j = 0; j < 4; j++) begin
            a[j]    = out[substage][j+subsubstage*4+0*16];
            b[j]    = out[substage][j+subsubstage*4+1*16];
            c[j]    = out[substage][j+subsubstage*4+2*16];
            d[j]    = out[substage][j+subsubstage*4+3*16];
            w0[j]   = w_256[substage*(j+subsubstage*4+0*16)];
            w1[j]   = w_256[substage*(j+subsubstage*4+1*16)];
            w2[j]   = w_256[substage*(j+subsubstage*4+2*16)];
            w3[j]   = w_256[substage*(j+subsubstage*4+3*16)];
        end
    end

    STAGE3: begin
        // for (int i = 0; i < 4; i++) begin
        //     for (int j = 0; j < 4; j++) begin
        //         for (int k = 0; k < 4; k++) begin
        //             a[i*16+j*4+k] = out[j][i*16+k+0*4];
        //             b[i*16+j*4+k] = out[j][i*16+k+1*4];
        //             c[i*16+j*4+k] = out[j][i*16+k+2*4];
        //             d[i*16+j*4+k] = out[j][i*16+k+3*4];
        //             w0[i*16+j*4+k]= w_256[j*4*(k+0*4)];
        //             w1[i*16+j*4+k]= w_256[j*4*(k+1*4)];
        //             w2[i*16+j*4+k]= w_256[j*4*(k+2*4)];
        //             w3[i*16+j*4+k]= w_256[j*4*(k+3*4)];
        //         end
        //     end
        // end
        for (int k = 0; k < 4; k++) begin
            a[k]    = out[subsubstage][substage*16+k+0*4];
            b[k]    = out[subsubstage][substage*16+k+1*4];
            c[k]    = out[subsubstage][substage*16+k+2*4];
            d[k]    = out[subsubstage][substage*16+k+3*4];
            w0[k]   = w_256[subsubstage*4*(k+0*4)];
            w1[k]   = w_256[subsubstage*4*(k+1*4)];
            w2[k]   = w_256[subsubstage*4*(k+2*4)];
            w3[k]   = w_256[subsubstage*4*(k+3*4)];
        end
    end

    STAGE4: begin
        // for (int i = 0; i < 4; i++) begin
        //     for (int j = 0; j < 4; j++) begin
        //         for (int k = 0; k < 4; k++) begin
        //             a[i*16+j*4+k] = out[k][i*16+j*4+0];
        //             b[i*16+j*4+k] = out[k][i*16+j*4+1];
        //             c[i*16+j*4+k] = out[k][i*16+j*4+2];
        //             d[i*16+j*4+k] = out[k][i*16+j*4+3];
        //             w0[i*16+j*4+k]= w_256[k*0*16];
        //             w1[i*16+j*4+k]= w_256[k*1*16];
        //             w2[i*16+j*4+k]= w_256[k*2*16];
        //             w3[i*16+j*4+k]= w_256[k*3*16];
        //         end
        //     end
        // end
        for (int k = 0; k < 4; k++) begin
            a[k]    = out[k][substage*16+subsubstage*4+0];
            b[k]    = out[k][substage*16+subsubstage*4+1];
            c[k]    = out[k][substage*16+subsubstage*4+2];
            d[k]    = out[k][substage*16+subsubstage*4+3];
            w0[k]   = w_256[k*0*16];
            w1[k]   = w_256[k*1*16];
            w2[k]   = w_256[k*2*16];
            w3[k]   = w_256[k*3*16];
        end
    end

    DONE: begin
        for (int i = 0; i < N_INST; i++) begin
            a[i] = 1'b0;
            b[i] = 1'b0;
            c[i] = 1'b0;
            d[i] = 1'b0;
            w0[i]= 1'b0;
            w1[i]= 1'b0;
            w2[i]= 1'b0;
            w3[i]= 1'b0;
        end
    end

    default: begin
        for (int i = 0; i < N_INST; i++) begin
            a[i] = 1'b0;
            b[i] = 1'b0;
            c[i] = 1'b0;
            d[i] = 1'b0;
            w0[i]= 1'b0;
            w1[i]= 1'b0;
            w2[i]= 1'b0;
            w3[i]= 1'b0;
        end

    end
    endcase
end

// state transition logic 
always_comb begin
    case (state)
    SET: begin
        if (start) begin
            state_d = STAGE1;
        end else begin
            state_d = SET;
        end
    end

    STAGE1: begin
        if (rst) begin
            state_d = SET;  
        end else if (counter == 4'hf) begin
            state_d = STAGE2;
        end else begin
            state_d = STAGE1;
        end
    end

    STAGE2: begin
        if (rst) begin
            state_d = SET;
        end else if (counter == 4'hf) begin
            state_d = STAGE3;
        end else begin 
            state_d = STAGE2;
        end
    end

    STAGE3: begin
        if (rst) begin
            state_d = SET;
        end else if (counter == 4'hf) begin 
            state_d = STAGE4;
        end else begin
            state_d = STAGE3;
        end
    end

    STAGE4: begin
        if (rst) begin 
            state_d = SET;
        end else if (counter == 4'hf) begin
            state_d = DONE;
        end else begin
            state_d = STAGE4;
        end
    end

    DONE: begin
        // if (rst) begin
        //     state_d = SET;
        // end else begin
        //     state_d = DONE;
        // end
        if (counter == 4'hf) begin
            state_d = SET;
        end else begin
            state_d = DONE;
        end
    end

    default: begin
        state_d = SET;
    end

    endcase
end

// catch frequency outputs
always_ff @(negedge clk) begin
    if (done_sr == 2'b10) begin
        for (int i = 0; i < 4; i++) begin
            for (int j = 0; j < 4; j++) begin
                for (int k = 0; k < 4; k++) begin
                    freq_real[i+j*4+k*16+N_BFLY*0] <= out[0][i*16+j*4+k][FULL_WIDTH-1:WIDTH];
                    freq_real[i+j*4+k*16+N_BFLY*1] <= out[1][i*16+j*4+k][FULL_WIDTH-1:WIDTH];
                    freq_real[i+j*4+k*16+N_BFLY*2] <= out[2][i*16+j*4+k][FULL_WIDTH-1:WIDTH];
                    freq_real[i+j*4+k*16+N_BFLY*3] <= out[3][i*16+j*4+k][FULL_WIDTH-1:WIDTH];

                    freq_imag[i+j*4+k*16+N_BFLY*0] <= out[0][i*16+j*4+k][WIDTH-1:0];
                    freq_imag[i+j*4+k*16+N_BFLY*1] <= out[1][i*16+j*4+k][WIDTH-1:0];
                    freq_imag[i+j*4+k*16+N_BFLY*2] <= out[2][i*16+j*4+k][WIDTH-1:0];
                    freq_imag[i+j*4+k*16+N_BFLY*3] <= out[3][i*16+j*4+k][WIDTH-1:0];
                end
            end
        end
    end else if (rst) begin
        for (int i = 0; i < N; i++) begin
            freq_real[i] <= 1'b0;
            freq_imag[i] <= 1'b0;
        end
    end
end

endmodule